module riscv


