module main

fn main() {
	a := 0b1111111
	println(a)
	println('Hello World!')
}
