module riscv